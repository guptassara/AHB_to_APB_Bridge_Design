module AHB_Master (
    Hclk,
    Hresetn,
    Hresp,
    Hrdata,
    Hwrite,
    Hreadyin,
    Hreadyout,
    Htrans,
    Hwdata,
    Haddr
);

  input Hclk, Hresetn, Hreadyout;
  input [1:0] Hresp;
  input [31:0] Hrdata;
  output reg Hwrite, Hreadyin;
  output reg [1:0] Htrans;
  output reg [31:0] Hwdata, Haddr;

  reg [2:0] Hburst;
  reg [2:0] Hsize;



  task single_write();
    begin
      @(posedge Hclk) #2;
      begin
        Hwrite = 1;
        Htrans = 2'b10;
        Hsize = 3'b000;
        Hburst = 3'b000;
        Hreadyin = 1;
        Haddr = 32'h8000_0001;
      end

      @(posedge Hclk) #2;
      begin
        Htrans = ($random)%256;
        Hwdata = ($random)%256;
      end
    end
  endtask


  task single_read();
    begin
      @(posedge Hclk) #2;
      begin
        Hwrite = 0;
        Htrans = 2'b10;
        Hsize = 3'b000;
        Hburst = 3'b000;
        Hreadyin = 1;
        Haddr = 32'h8000_00A2;
      end

      @(posedge Hclk) #2;
      begin
        Htrans = 2'b00;
      end
    end
  endtask


endmodule
